magic
tech scmos
timestamp 1593967954
<< metal1 >>
rect 99 89 103 90
rect 99 85 111 89
rect 99 81 103 85
rect 60 77 103 81
rect 60 75 64 77
rect -16 39 0 43
rect 102 40 106 62
rect -16 6 -12 39
rect 95 36 106 40
rect 177 39 181 41
rect 95 16 98 36
rect 60 13 98 16
rect 101 6 106 13
rect -18 2 -12 6
rect 60 4 106 6
rect 64 2 106 4
rect -16 -31 -12 2
rect -16 -35 -4 -31
rect 102 -34 106 -21
rect 96 -37 107 -34
rect 96 -55 99 -37
rect 64 -59 99 -55
rect 102 -68 107 -60
rect 181 -65 186 -62
<< m2contact >>
rect 95 43 99 48
rect 95 -31 99 -26
rect 151 -30 159 -24
rect 214 -28 219 -24
<< metal2 >>
rect 99 44 219 47
rect 215 -24 219 44
rect 99 -30 151 -26
use vsdswitch  vsdswitch_0
timestamp 1593965765
transform 1 0 10 0 1 47
box -17 -32 89 32
use resistor2  resistor2_0
timestamp 1593964240
transform 1 0 114 0 1 79
box -9 -22 36 11
use resistor2  resistor2_1
timestamp 1593964240
transform 1 0 109 0 1 30
box -9 -22 36 11
use vsdswitch  vsdswitch_1
timestamp 1593965765
transform 1 0 10 0 1 -27
box -17 -32 89 32
use resistor2  resistor2_2
timestamp 1593964240
transform 1 0 110 0 1 -4
box -9 -22 36 11
use resistor2  resistor2_3
timestamp 1593964240
transform 1 0 110 0 1 -43
box -9 -22 36 11
use vsdswitch  vsdswitch_2
timestamp 1593965765
transform 0 1 185 -1 0 26
box -17 -32 89 32
<< labels >>
rlabel metal1 -18 2 -18 6 3 D0!
rlabel metal1 102 -68 107 -68 1 res_out
rlabel metal1 99 90 103 90 5 res_in
rlabel metal1 177 41 181 41 1 D1!
rlabel metal1 181 -65 186 -65 1 output
<< end >>
