* SPICE3 file created from 5bitres.ext - technology: scmos

.option scale=0.1u

R0 4bitres_1/3bitres_0/2bitres_0/resistor2_1/a 4bitres_1/3bitres_0/2bitres_0/res_in polyResistor w=2 l=263
R1 4bitres_1/3bitres_0/2bitres_0/resistor2_1/b 4bitres_1/3bitres_0/2bitres_0/resistor2_1/a polyResistor w=2 l=263
M1000 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/in_1 4bitres_1/3bitres_0/2bitres_0/vsdswitch_0/invout 4bitres_1/3bitres_0/2bitres_0/resistor2_1/a gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 4bitres_1/3bitres_0/2bitres_0/res_in D0 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 4bitres_1/3bitres_0/2bitres_0/resistor2_1/a D0 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/in_1 4bitres_1/3bitres_0/2bitres_0/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 4bitres_1/3bitres_0/2bitres_0/vsdswitch_0/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 4bitres_1/3bitres_0/2bitres_0/vsdswitch_0/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/in_1 4bitres_1/3bitres_0/2bitres_0/vsdswitch_0/invout 4bitres_1/3bitres_0/2bitres_0/res_in 4bitres_1/3bitres_0/2bitres_0/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R2 4bitres_1/3bitres_0/2bitres_1/res_in 4bitres_1/3bitres_0/2bitres_0/resistor2_2/b polyResistor w=2 l=263
R3 4bitres_1/3bitres_0/2bitres_0/resistor2_2/b 4bitres_1/3bitres_0/2bitres_0/resistor2_1/b polyResistor w=2 l=263
M1006 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/VOUT 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/invout 4bitres_1/3bitres_0/2bitres_0/resistor2_2/b gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 4bitres_1/3bitres_0/2bitres_0/resistor2_1/b D0 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 4bitres_1/3bitres_0/2bitres_0/resistor2_2/b D0 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/VOUT 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/VOUT 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/invout 4bitres_1/3bitres_0/2bitres_0/resistor2_1/b 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 4bitres_1/3bitres_0/2bitres_0/output 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/invout 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/in_1 D1 4bitres_1/3bitres_0/2bitres_0/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 4bitres_1/3bitres_0/2bitres_0/vsdswitch_1/VOUT D1 4bitres_1/3bitres_0/2bitres_0/output 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/invout D1 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/invout D1 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 4bitres_1/3bitres_0/2bitres_0/output 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/invout 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/in_1 4bitres_1/3bitres_0/2bitres_0/vsdswitch_2/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R4 4bitres_1/3bitres_0/2bitres_1/resistor2_1/a 4bitres_1/3bitres_0/2bitres_1/res_in polyResistor w=2 l=263
R5 4bitres_1/3bitres_0/2bitres_1/resistor2_1/b 4bitres_1/3bitres_0/2bitres_1/resistor2_1/a polyResistor w=2 l=263
M1018 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/in_1 4bitres_1/3bitres_0/2bitres_1/vsdswitch_0/invout 4bitres_1/3bitres_0/2bitres_1/resistor2_1/a gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 4bitres_1/3bitres_0/2bitres_1/res_in D0 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 4bitres_1/3bitres_0/2bitres_1/resistor2_1/a D0 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/in_1 4bitres_1/3bitres_0/2bitres_1/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 4bitres_1/3bitres_0/2bitres_1/vsdswitch_0/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 4bitres_1/3bitres_0/2bitres_1/vsdswitch_0/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/in_1 4bitres_1/3bitres_0/2bitres_1/vsdswitch_0/invout 4bitres_1/3bitres_0/2bitres_1/res_in 4bitres_1/3bitres_0/2bitres_1/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R6 4bitres_1/3bitres_1/2bitres_0/res_in 4bitres_1/3bitres_0/2bitres_1/resistor2_2/b polyResistor w=2 l=263
R7 4bitres_1/3bitres_0/2bitres_1/resistor2_2/b 4bitres_1/3bitres_0/2bitres_1/resistor2_1/b polyResistor w=2 l=263
M1024 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/VOUT 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/invout 4bitres_1/3bitres_0/2bitres_1/resistor2_2/b gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 4bitres_1/3bitres_0/2bitres_1/resistor2_1/b D0 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 4bitres_1/3bitres_0/2bitres_1/resistor2_2/b D0 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/VOUT 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1029 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/VOUT 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/invout 4bitres_1/3bitres_0/2bitres_1/resistor2_1/b 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 4bitres_1/3bitres_0/2bitres_1/output 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/invout 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/in_1 D1 4bitres_1/3bitres_0/2bitres_1/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 4bitres_1/3bitres_0/2bitres_1/vsdswitch_1/VOUT D1 4bitres_1/3bitres_0/2bitres_1/output 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1033 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/invout D1 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/invout D1 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1035 4bitres_1/3bitres_0/2bitres_1/output 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/invout 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/in_1 4bitres_1/3bitres_0/2bitres_1/vsdswitch_2/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 4bitres_1/vsdswitch_0/in_1 4bitres_1/3bitres_0/vsdswitch_0/invout 4bitres_1/3bitres_0/2bitres_1/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 4bitres_1/3bitres_0/2bitres_0/output D2 4bitres_1/vsdswitch_0/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 4bitres_1/3bitres_0/2bitres_1/output D2 4bitres_1/vsdswitch_0/in_1 4bitres_1/3bitres_0/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 4bitres_1/3bitres_0/vsdswitch_0/invout D2 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 4bitres_1/3bitres_0/vsdswitch_0/invout D2 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 4bitres_1/vsdswitch_0/in_1 4bitres_1/3bitres_0/vsdswitch_0/invout 4bitres_1/3bitres_0/2bitres_0/output 4bitres_1/3bitres_0/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R8 4bitres_1/3bitres_1/2bitres_0/resistor2_1/a 4bitres_1/3bitres_1/2bitres_0/res_in polyResistor w=2 l=263
R9 4bitres_1/3bitres_1/2bitres_0/resistor2_1/b 4bitres_1/3bitres_1/2bitres_0/resistor2_1/a polyResistor w=2 l=263
M1042 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/in_1 4bitres_1/3bitres_1/2bitres_0/vsdswitch_0/invout 4bitres_1/3bitres_1/2bitres_0/resistor2_1/a gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 4bitres_1/3bitres_1/2bitres_0/res_in D0 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 4bitres_1/3bitres_1/2bitres_0/resistor2_1/a D0 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/in_1 4bitres_1/3bitres_1/2bitres_0/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 4bitres_1/3bitres_1/2bitres_0/vsdswitch_0/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 4bitres_1/3bitres_1/2bitres_0/vsdswitch_0/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1047 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/in_1 4bitres_1/3bitres_1/2bitres_0/vsdswitch_0/invout 4bitres_1/3bitres_1/2bitres_0/res_in 4bitres_1/3bitres_1/2bitres_0/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R10 4bitres_1/3bitres_1/2bitres_1/res_in 4bitres_1/3bitres_1/2bitres_0/resistor2_2/b polyResistor w=2 l=263
R11 4bitres_1/3bitres_1/2bitres_0/resistor2_2/b 4bitres_1/3bitres_1/2bitres_0/resistor2_1/b polyResistor w=2 l=263
M1048 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/VOUT 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/invout 4bitres_1/3bitres_1/2bitres_0/resistor2_2/b gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1049 4bitres_1/3bitres_1/2bitres_0/resistor2_1/b D0 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 4bitres_1/3bitres_1/2bitres_0/resistor2_2/b D0 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/VOUT 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/VOUT 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/invout 4bitres_1/3bitres_1/2bitres_0/resistor2_1/b 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 4bitres_1/3bitres_1/2bitres_0/output 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/invout 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/in_1 D1 4bitres_1/3bitres_1/2bitres_0/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 4bitres_1/3bitres_1/2bitres_0/vsdswitch_1/VOUT D1 4bitres_1/3bitres_1/2bitres_0/output 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1057 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/invout D1 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/invout D1 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1059 4bitres_1/3bitres_1/2bitres_0/output 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/invout 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/in_1 4bitres_1/3bitres_1/2bitres_0/vsdswitch_2/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R12 4bitres_1/3bitres_1/2bitres_1/resistor2_1/a 4bitres_1/3bitres_1/2bitres_1/res_in polyResistor w=2 l=263
R13 4bitres_1/3bitres_1/2bitres_1/resistor2_1/b 4bitres_1/3bitres_1/2bitres_1/resistor2_1/a polyResistor w=2 l=263
M1060 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/in_1 4bitres_1/3bitres_1/2bitres_1/vsdswitch_0/invout 4bitres_1/3bitres_1/2bitres_1/resistor2_1/a gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1061 4bitres_1/3bitres_1/2bitres_1/res_in D0 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 4bitres_1/3bitres_1/2bitres_1/resistor2_1/a D0 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/in_1 4bitres_1/3bitres_1/2bitres_1/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 4bitres_1/3bitres_1/2bitres_1/vsdswitch_0/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 4bitres_1/3bitres_1/2bitres_1/vsdswitch_0/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/in_1 4bitres_1/3bitres_1/2bitres_1/vsdswitch_0/invout 4bitres_1/3bitres_1/2bitres_1/res_in 4bitres_1/3bitres_1/2bitres_1/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R14 4bitres_1/3bitres_1/2bitres_1/res_out 4bitres_1/3bitres_1/2bitres_1/resistor2_2/b polyResistor w=2 l=263
R15 4bitres_1/3bitres_1/2bitres_1/resistor2_2/b 4bitres_1/3bitres_1/2bitres_1/resistor2_1/b polyResistor w=2 l=263
M1066 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/VOUT 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/invout 4bitres_1/3bitres_1/2bitres_1/resistor2_2/b gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 4bitres_1/3bitres_1/2bitres_1/resistor2_1/b D0 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 4bitres_1/3bitres_1/2bitres_1/resistor2_2/b D0 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/VOUT 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1071 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/VOUT 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/invout 4bitres_1/3bitres_1/2bitres_1/resistor2_1/b 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 4bitres_1/3bitres_1/2bitres_1/output 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/invout 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/in_1 D1 4bitres_1/3bitres_1/2bitres_1/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 4bitres_1/3bitres_1/2bitres_1/vsdswitch_1/VOUT D1 4bitres_1/3bitres_1/2bitres_1/output 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/invout D1 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/invout D1 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 4bitres_1/3bitres_1/2bitres_1/output 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/invout 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/in_1 4bitres_1/3bitres_1/2bitres_1/vsdswitch_2/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 4bitres_1/vsdswitch_0/in_2 4bitres_1/3bitres_1/vsdswitch_0/invout 4bitres_1/3bitres_1/2bitres_1/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 4bitres_1/3bitres_1/2bitres_0/output D2 4bitres_1/vsdswitch_0/in_2 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 4bitres_1/3bitres_1/2bitres_1/output D2 4bitres_1/vsdswitch_0/in_2 4bitres_1/3bitres_1/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 4bitres_1/3bitres_1/vsdswitch_0/invout D2 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 4bitres_1/3bitres_1/vsdswitch_0/invout D2 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 4bitres_1/vsdswitch_0/in_2 4bitres_1/3bitres_1/vsdswitch_0/invout 4bitres_1/3bitres_1/2bitres_0/output 4bitres_1/3bitres_1/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1084 vsdswitch_0/in_2 4bitres_1/vsdswitch_0/invout 4bitres_1/vsdswitch_0/in_2 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 4bitres_1/vsdswitch_0/in_1 D3 vsdswitch_0/in_2 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 4bitres_1/vsdswitch_0/in_2 D3 vsdswitch_0/in_2 4bitres_1/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 4bitres_1/vsdswitch_0/invout D3 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 4bitres_1/vsdswitch_0/invout D3 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 vsdswitch_0/in_2 4bitres_1/vsdswitch_0/invout 4bitres_1/vsdswitch_0/in_1 4bitres_1/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 out_five vsdswitch_0/invout vsdswitch_0/in_2 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 vsdswitch_0/in_1 D4 out_five gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1092 vsdswitch_0/in_2 D4 out_five vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1093 vsdswitch_0/invout D4 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 vsdswitch_0/invout D4 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 out_five vsdswitch_0/invout vsdswitch_0/in_1 vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R16 4bitres_0/3bitres_0/2bitres_0/resistor2_1/a 4bitres_0/3bitres_0/2bitres_0/res_in polyResistor w=2 l=263
R17 4bitres_0/3bitres_0/2bitres_0/resistor2_1/b 4bitres_0/3bitres_0/2bitres_0/resistor2_1/a polyResistor w=2 l=263
M1096 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/in_1 4bitres_0/3bitres_0/2bitres_0/vsdswitch_0/invout 4bitres_0/3bitres_0/2bitres_0/resistor2_1/a gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1097 4bitres_0/3bitres_0/2bitres_0/res_in D0 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1098 4bitres_0/3bitres_0/2bitres_0/resistor2_1/a D0 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/in_1 4bitres_0/3bitres_0/2bitres_0/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 4bitres_0/3bitres_0/2bitres_0/vsdswitch_0/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 4bitres_0/3bitres_0/2bitres_0/vsdswitch_0/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/in_1 4bitres_0/3bitres_0/2bitres_0/vsdswitch_0/invout 4bitres_0/3bitres_0/2bitres_0/res_in 4bitres_0/3bitres_0/2bitres_0/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R18 4bitres_0/3bitres_0/2bitres_1/res_in 4bitres_0/3bitres_0/2bitres_0/resistor2_2/b polyResistor w=2 l=263
R19 4bitres_0/3bitres_0/2bitres_0/resistor2_2/b 4bitres_0/3bitres_0/2bitres_0/resistor2_1/b polyResistor w=2 l=263
M1102 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/VOUT 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/invout 4bitres_0/3bitres_0/2bitres_0/resistor2_2/b gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 4bitres_0/3bitres_0/2bitres_0/resistor2_1/b D0 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 4bitres_0/3bitres_0/2bitres_0/resistor2_2/b D0 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/VOUT 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1105 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1107 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/VOUT 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/invout 4bitres_0/3bitres_0/2bitres_0/resistor2_1/b 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 4bitres_0/3bitres_0/2bitres_0/output 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/invout 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/in_1 D1 4bitres_0/3bitres_0/2bitres_0/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 4bitres_0/3bitres_0/2bitres_0/vsdswitch_1/VOUT D1 4bitres_0/3bitres_0/2bitres_0/output 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/invout D1 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/invout D1 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 4bitres_0/3bitres_0/2bitres_0/output 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/invout 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/in_1 4bitres_0/3bitres_0/2bitres_0/vsdswitch_2/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R20 4bitres_0/3bitres_0/2bitres_1/resistor2_1/a 4bitres_0/3bitres_0/2bitres_1/res_in polyResistor w=2 l=263
R21 4bitres_0/3bitres_0/2bitres_1/resistor2_1/b 4bitres_0/3bitres_0/2bitres_1/resistor2_1/a polyResistor w=2 l=263
M1114 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/in_1 4bitres_0/3bitres_0/2bitres_1/vsdswitch_0/invout 4bitres_0/3bitres_0/2bitres_1/resistor2_1/a gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 4bitres_0/3bitres_0/2bitres_1/res_in D0 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 4bitres_0/3bitres_0/2bitres_1/resistor2_1/a D0 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/in_1 4bitres_0/3bitres_0/2bitres_1/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1117 4bitres_0/3bitres_0/2bitres_1/vsdswitch_0/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 4bitres_0/3bitres_0/2bitres_1/vsdswitch_0/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/in_1 4bitres_0/3bitres_0/2bitres_1/vsdswitch_0/invout 4bitres_0/3bitres_0/2bitres_1/res_in 4bitres_0/3bitres_0/2bitres_1/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R22 4bitres_0/3bitres_1/2bitres_0/res_in 4bitres_0/3bitres_0/2bitres_1/resistor2_2/b polyResistor w=2 l=263
R23 4bitres_0/3bitres_0/2bitres_1/resistor2_2/b 4bitres_0/3bitres_0/2bitres_1/resistor2_1/b polyResistor w=2 l=263
M1120 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/VOUT 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/invout 4bitres_0/3bitres_0/2bitres_1/resistor2_2/b gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 4bitres_0/3bitres_0/2bitres_1/resistor2_1/b D0 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 4bitres_0/3bitres_0/2bitres_1/resistor2_2/b D0 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/VOUT 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/VOUT 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/invout 4bitres_0/3bitres_0/2bitres_1/resistor2_1/b 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1126 4bitres_0/3bitres_0/2bitres_1/output 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/invout 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/in_1 D1 4bitres_0/3bitres_0/2bitres_1/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 4bitres_0/3bitres_0/2bitres_1/vsdswitch_1/VOUT D1 4bitres_0/3bitres_0/2bitres_1/output 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/invout D1 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/invout D1 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 4bitres_0/3bitres_0/2bitres_1/output 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/invout 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/in_1 4bitres_0/3bitres_0/2bitres_1/vsdswitch_2/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 4bitres_0/vsdswitch_0/in_1 4bitres_0/3bitres_0/vsdswitch_0/invout 4bitres_0/3bitres_0/2bitres_1/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 4bitres_0/3bitres_0/2bitres_0/output D2 4bitres_0/vsdswitch_0/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 4bitres_0/3bitres_0/2bitres_1/output D2 4bitres_0/vsdswitch_0/in_1 4bitres_0/3bitres_0/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 4bitres_0/3bitres_0/vsdswitch_0/invout D2 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 4bitres_0/3bitres_0/vsdswitch_0/invout D2 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1137 4bitres_0/vsdswitch_0/in_1 4bitres_0/3bitres_0/vsdswitch_0/invout 4bitres_0/3bitres_0/2bitres_0/output 4bitres_0/3bitres_0/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R24 4bitres_0/3bitres_1/2bitres_0/resistor2_1/a 4bitres_0/3bitres_1/2bitres_0/res_in polyResistor w=2 l=263
R25 4bitres_0/3bitres_1/2bitres_0/resistor2_1/b 4bitres_0/3bitres_1/2bitres_0/resistor2_1/a polyResistor w=2 l=263
M1138 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/in_1 4bitres_0/3bitres_1/2bitres_0/vsdswitch_0/invout 4bitres_0/3bitres_1/2bitres_0/resistor2_1/a gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 4bitres_0/3bitres_1/2bitres_0/res_in D0 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 4bitres_0/3bitres_1/2bitres_0/resistor2_1/a D0 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/in_1 4bitres_0/3bitres_1/2bitres_0/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 4bitres_0/3bitres_1/2bitres_0/vsdswitch_0/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 4bitres_0/3bitres_1/2bitres_0/vsdswitch_0/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1143 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/in_1 4bitres_0/3bitres_1/2bitres_0/vsdswitch_0/invout 4bitres_0/3bitres_1/2bitres_0/res_in 4bitres_0/3bitres_1/2bitres_0/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R26 4bitres_0/3bitres_1/2bitres_1/res_in 4bitres_0/3bitres_1/2bitres_0/resistor2_2/b polyResistor w=2 l=263
R27 4bitres_0/3bitres_1/2bitres_0/resistor2_2/b 4bitres_0/3bitres_1/2bitres_0/resistor2_1/b polyResistor w=2 l=263
M1144 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/VOUT 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/invout 4bitres_0/3bitres_1/2bitres_0/resistor2_2/b gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 4bitres_0/3bitres_1/2bitres_0/resistor2_1/b D0 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 4bitres_0/3bitres_1/2bitres_0/resistor2_2/b D0 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/VOUT 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1149 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/VOUT 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/invout 4bitres_0/3bitres_1/2bitres_0/resistor2_1/b 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 4bitres_0/3bitres_1/2bitres_0/output 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/invout 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1151 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/in_1 D1 4bitres_0/3bitres_1/2bitres_0/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 4bitres_0/3bitres_1/2bitres_0/vsdswitch_1/VOUT D1 4bitres_0/3bitres_1/2bitres_0/output 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/invout D1 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/invout D1 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 4bitres_0/3bitres_1/2bitres_0/output 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/invout 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/in_1 4bitres_0/3bitres_1/2bitres_0/vsdswitch_2/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R28 4bitres_0/3bitres_1/2bitres_1/resistor2_1/a 4bitres_0/3bitres_1/2bitres_1/res_in polyResistor w=2 l=263
R29 4bitres_0/3bitres_1/2bitres_1/resistor2_1/b 4bitres_0/3bitres_1/2bitres_1/resistor2_1/a polyResistor w=2 l=263
M1156 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/in_1 4bitres_0/3bitres_1/2bitres_1/vsdswitch_0/invout 4bitres_0/3bitres_1/2bitres_1/resistor2_1/a gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1157 4bitres_0/3bitres_1/2bitres_1/res_in D0 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 4bitres_0/3bitres_1/2bitres_1/resistor2_1/a D0 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/in_1 4bitres_0/3bitres_1/2bitres_1/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 4bitres_0/3bitres_1/2bitres_1/vsdswitch_0/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 4bitres_0/3bitres_1/2bitres_1/vsdswitch_0/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1161 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/in_1 4bitres_0/3bitres_1/2bitres_1/vsdswitch_0/invout 4bitres_0/3bitres_1/2bitres_1/res_in 4bitres_0/3bitres_1/2bitres_1/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
R30 4bitres_1/3bitres_0/2bitres_0/res_in 4bitres_0/3bitres_1/2bitres_1/resistor2_2/b polyResistor w=2 l=263
R31 4bitres_0/3bitres_1/2bitres_1/resistor2_2/b 4bitres_0/3bitres_1/2bitres_1/resistor2_1/b polyResistor w=2 l=263
M1162 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/VOUT 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/invout 4bitres_0/3bitres_1/2bitres_1/resistor2_2/b gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1163 4bitres_0/3bitres_1/2bitres_1/resistor2_1/b D0 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 4bitres_0/3bitres_1/2bitres_1/resistor2_2/b D0 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/VOUT 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/invout D0 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/invout D0 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/VOUT 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/invout 4bitres_0/3bitres_1/2bitres_1/resistor2_1/b 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 4bitres_0/3bitres_1/2bitres_1/output 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/invout 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/VOUT gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1169 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/in_1 D1 4bitres_0/3bitres_1/2bitres_1/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 4bitres_0/3bitres_1/2bitres_1/vsdswitch_1/VOUT D1 4bitres_0/3bitres_1/2bitres_1/output 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/invout D1 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/invout D1 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 4bitres_0/3bitres_1/2bitres_1/output 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/invout 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/in_1 4bitres_0/3bitres_1/2bitres_1/vsdswitch_2/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 4bitres_0/vsdswitch_0/in_2 4bitres_0/3bitres_1/vsdswitch_0/invout 4bitres_0/3bitres_1/2bitres_1/output gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 4bitres_0/3bitres_1/2bitres_0/output D2 4bitres_0/vsdswitch_0/in_2 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 4bitres_0/3bitres_1/2bitres_1/output D2 4bitres_0/vsdswitch_0/in_2 4bitres_0/3bitres_1/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 4bitres_0/3bitres_1/vsdswitch_0/invout D2 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 4bitres_0/3bitres_1/vsdswitch_0/invout D2 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 4bitres_0/vsdswitch_0/in_2 4bitres_0/3bitres_1/vsdswitch_0/invout 4bitres_0/3bitres_1/2bitres_0/output 4bitres_0/3bitres_1/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1180 vsdswitch_0/in_1 4bitres_0/vsdswitch_0/invout 4bitres_0/vsdswitch_0/in_2 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 4bitres_0/vsdswitch_0/in_1 D3 vsdswitch_0/in_1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 4bitres_0/vsdswitch_0/in_2 D3 vsdswitch_0/in_1 4bitres_0/vsdswitch_0/w_57_n21# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 4bitres_0/vsdswitch_0/invout D3 vdd vdd pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1184 4bitres_0/vsdswitch_0/invout D3 gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 vsdswitch_0/in_1 4bitres_0/vsdswitch_0/invout 4bitres_0/vsdswitch_0/in_1 4bitres_0/vsdswitch_0/w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
