* SPICE3 file created from vsdswitch.ext - technology: scmos

.option scale=0.1u

M1000 VOUT invout in_2 gnd nfet w=4 l=2
+  ad=56 pd=44 as=28 ps=22
M1001 in_1 dig_in VOUT gnd nfet w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1002 in_2 dig_in VOUT w_57_n21# pfet w=9 l=2
+  ad=63 pd=32 as=126 ps=64
M1003 invout dig_in vdd vdd pfet w=9 l=2
+  ad=63 pd=32 as=63 ps=32
M1004 invout dig_in gnd gnd nfet w=4 l=2
+  ad=28 pd=22 as=28 ps=22
M1005 VOUT invout in_1 w_21_1# pfet w=9 l=2
+  ad=0 pd=0 as=63 ps=32
