magic
tech scmos
timestamp 1593964240
<< polycontact >>
rect -8 6 -3 10
rect -8 -21 -3 -17
<< pseudo_rpoly >>
rect -9 10 36 11
rect -9 6 -8 10
rect -3 8 36 10
rect -9 5 33 6
rect -9 4 21 5
rect 23 4 33 5
rect -9 3 33 4
rect -9 -4 -8 3
rect 35 1 36 8
rect -6 -2 36 1
rect -9 -5 33 -4
rect -9 -6 21 -5
rect 23 -6 33 -5
rect -9 -7 33 -6
rect -9 -14 -8 -7
rect 35 -9 36 -2
rect -6 -12 36 -9
rect -9 -15 33 -14
rect -9 -16 21 -15
rect 23 -16 33 -15
rect -9 -17 33 -16
rect -9 -21 -8 -17
rect 35 -19 36 -12
rect -3 -21 36 -19
rect -9 -22 36 -21
<< rpoly >>
rect -3 6 35 8
rect 33 3 35 6
rect -8 1 35 3
rect -8 -2 -6 1
rect -8 -4 35 -2
rect 33 -7 35 -4
rect -8 -9 35 -7
rect -8 -12 -6 -9
rect -8 -14 35 -12
rect 33 -17 35 -14
rect -3 -19 35 -17
<< labels >>
rlabel polycontact -6 8 -6 8 4 a
rlabel polycontact -5 -19 -5 -19 2 b
<< end >>
